library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity RF_DestReg_Decoder_20332706 is
    Port ( 
        A : in std_logic_vector(4 downto 0);
        D : out std_logic_vector(31 downto 0)
   );
end RF_DestReg_Decoder_20332706;

architecture Behavioral of RF_DestReg_Decoder_20332706 is
    begin
        process(A)
        begin
            case A is
                WHEN "00000" => D <= "00000000000000000000000000000001";
                WHEN "00001" => D <= "00000000000000000000000000000010";
                WHEN "00010" => D <= "00000000000000000000000000000100";
                WHEN "00011" => D <= "00000000000000000000000000001000";
                WHEN "00100" => D <= "00000000000000000000000000010000";
                WHEN "00101" => D <= "00000000000000000000000000100000";
                WHEN "00110" => D <= "00000000000000000000000001000000";
                WHEN "00111" => D <= "00000000000000000000000010000000";
                WHEN "01000" => D <= "00000000000000000000000100000000";
                WHEN "01001" => D <= "00000000000000000000001000000000";
                WHEN "01010" => D <= "00000000000000000000010000000000";
                WHEN "01011" => D <= "00000000000000000000100000000000";
                WHEN "01100" => D <= "00000000000000000001000000000000";
                WHEN "01101" => D <= "00000000000000000010000000000000";
                WHEN "01110" => D <= "00000000000000000100000000000000";
                WHEN "01111" => D <= "00000000000000001000000000000000";
                WHEN "10000" => D <= "00000000000000010000000000000000";
                WHEN "10001" => D <= "00000000000000100000000000000000";
                WHEN "10010" => D <= "00000000000001000000000000000000";
                WHEN "10011" => D <= "00000000000010000000000000000000";
                WHEN "10100" => D <= "00000000000100000000000000000000";
                WHEN "10101" => D <= "00000000001000000000000000000000";
                WHEN "10110" => D <= "00000000010000000000000000000000";
                WHEN "10111" => D <= "00000000100000000000000000000000";
                WHEN "11000" => D <= "00000001000000000000000000000000";
                WHEN "11001" => D <= "00000010000000000000000000000000";
                WHEN "11010" => D <= "00000100000000000000000000000000";
                WHEN "11011" => D <= "00001000000000000000000000000000";
                WHEN "11100" => D <= "00010000000000000000000000000000";
                WHEN "11101" => D <= "00100000000000000000000000000000";
                WHEN "11110" => D <= "01000000000000000000000000000000";
                WHEN "11111" => D <= "10000000000000000000000000000000";
                WHEN OTHERS  => D <= "00000000000000000000000000000000";
            end case;
        end process;
end Behavioral;